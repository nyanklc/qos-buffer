module DisplayM(clock_50, clock_25, in_number, received1, received2, 
                received3, received4, dropped1, dropped2, dropped3, 
                dropped4, data1, data2, data3, data4, output_count1, output_count2, output_count3, output_count4, 
					 outputted_buffer_packet, red_sig, green_sig, blue_sig, hsync, vsync, nsync);
					 
	input clock_50;
	input clock_25;
	input wire[3:0] in_number;
	input wire[11:0] received1;
	input wire[11:0] received2;
	input wire[11:0] received3;
	input wire[11:0] received4;
	input wire[11:0] dropped1;
	input wire[11:0] dropped2;
	input wire[11:0] dropped3;
	input wire[11:0] dropped4;
	input wire[17:0] data1;
	input wire[17:0] data2;
	input wire[17:0] data3;
	input wire[17:0] data4;
	input wire[11:0] output_count1;
	input wire[11:0] output_count2;
	input wire[11:0] output_count3;
	input wire[11:0] output_count4;
	input wire[3:0] outputted_buffer_packet;
	 
	output red_sig;
	output green_sig;
	output blue_sig;
	
	reg red = 1;
	reg green = 1;
	reg blue = 1;
	 
	output hsync;
	output vsync;
	output nsync;
	 
	wire[15:0] hcount;
	wire[15:0] vcount;
	
	integer int_output_count1 = 0;
	integer int_output_count2 = 0;
	integer int_output_count3 = 0;
	integer int_output_count4 = 0;
	integer int_output_count_total = 0;
	integer int_received_count1 = 0;
	integer int_received_count2 = 0;
	integer int_received_count3 = 0;
	integer int_received_count4 = 0;
	integer int_received_count_total = 0;
	integer int_dropped_count1 = 0;
	integer int_dropped_count2 = 0;
	integer int_dropped_count3 = 0;
	integer int_dropped_count4 = 0;
	integer int_dropped_count_total = 0;
	integer dumdig = 0;
	
	reg[1599:0]block_sifir = 1600'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111110000000001111111111111111111111111111110000000000011111111111111111111111111110000011100001111111111111111111111111111000011110000011111111111111111111111111000011111100001111111111111111111111111100001111110000111111111111111111111111110000111111000011111111111111111111111111000011111100001111111111111111111111111100001111110000111111111111111111111111110000111111000011111111111111111111111111000011111100001111111111111111111111111100001111110000111111111111111111111111110000111111000011111111111111111111111111000011111100001111111111111111111111111100000111100000111111111111111111111111111000011110000111111111111111111111111111100000000000111111111111111111111111111111000000000011111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[1599:0]block_bir = 1600'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111100000011111111111111111111111111111111100000001111111111111111111111111111111100000000111111111111111111111111111111100001000011111111111111111111111111111110011100001111111111111111111111111111111111110000111111111111111111111111111111111111000011111111111111111111111111111111111100001111111111111111111111111111111111110000111111111111111111111111111111111111000011111111111111111111111111111111111100001111111111111111111111111111111111110000111111111111111111111111111111111111000011111111111111111111111111111111111100001111111111111111111111111111111111110000111111111111111111111111111111111111000011111111111111111111111111111111000000000000111111111111111111111111111100000000000011111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[1599:0]block_iki = 1600'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111100000000001111111111111111111111111111100000000000111111111111111111111111111110011110000001111111111111111111111111111011111100000111111111111111111111111111111111110000011111111111111111111111111111111111000001111111111111111111111111111111111100000111111111111111111111111111111111110000111111111111111111111111111111111110000011111111111111111111111111111111110000011111111111111111111111111111111111000001111111111111111111111111111111111000001111111111111111111111111111111111000001111111111111111111111111111111111000001111111111111111111111111111111111000001111111111111111111111111111111111000001111111111111111111111111111111111000000000000001111111111111111111111111100000000000000111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[1599:0]block_uc = 1600'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111100000000001111111111111111111111111111100000000000111111111111111111111111111110001111000001111111111111111111111111111011111100000111111111111111111111111111111111110000011111111111111111111111111111111111000001111111111111111111111111111111111000001111111111111111111111111111110000000001111111111111111111111111111111000000000111111111111111111111111111111100000000001111111111111111111111111111111111100000011111111111111111111111111111111111100000111111111111111111111111111111111110000011111111111111111111111111111111111000001111111111111111111111111111111111100000111111111111111111111111110011111100000111111111111111111111111111000000000000011111111111111111111111111100000000000011111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	
	reg[599:0]td_sifir = 600'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110000000011111111111100111100111111111110011111001111111111100111111001111111111001111110011111111110011111100111111111100111111001111111111001111110011111111110011111100111111111100111111001111111111001111100111111111111001111001111111111110001000111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[599:0]td_bir = 600'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111000111111111111111000001111111111111110010011111111111111111100111111111111111111001111111111111111110011111111111111111100111111111111111111001111111111111111110011111111111111111100111111111111111111001111111111111111110011111111111111111000011111111111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[599:0]td_iki = 600'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111100000001111111111111011110011111111111111111100011111111111111111000111111111111111110001111111111111111100111111111111111110001111111111111111100111111111111111110011111111111111111001111111111111111100111111111111111110011111111111111111000000000111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[599:0]td_uc = 600'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111100000001111111111111011110011111111111111111100011111111111111111000111111111111111110011111111111111000001111111111111110000011111111111111111110001111111111111111110011111111111111111100111111111111111111001111111111101111110011111111111000010001111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[599:0]td_dort = 600'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111100001111111111111111000011111111111111100100111111111111111001001111111111111100110011111111111111001100111111111111100111001111111111111011110011111111111100111100111111111111000100000111111111110000000000111111111111111100111111111111111111001111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[599:0]td_bes = 600'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111100000001111111111111001111111111111111110111111111111111111100111111111111111111000011111111111111110000000111111111111111111000111111111111111111001111111111111111110011111111111111111100111111111111111111001111111111111111100011111111111000000001111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[599:0]td_alti = 600'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111110000000111111111111000111111111111111110011111111111111111101111111111111111110011111111111111111100100000111111111111000000000111111111110011111000111111111100111111001111111111001111110011111111111011111100111111111110011110011111111111100000000111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[599:0]td_yedi = 600'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111111000000000011111111111111111001111111111111111110011111111111111111001111111111111111110011111111111111111001111111111111111110011111111111111111100111111111111111110011111111111111111100111111111111111110011111111111111111100111111111111111110001111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[599:0]td_sekiz = 600'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111100000000111111111111001111001111111111110111110011111111111100111100111111111111001110011111111111111000001111111111111111000011111111111111000100001111111111100011110011111111111001111110011111111110011111100111111111100111110011111111111100000000111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[599:0]td_dokuz = 600'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111110000000111111111111001111100111111111110011111001111111111100111110011111111111001111100011111111110011111000111111111110000000001111111111110000000111111111111111111001111111111111111110011111111111111111100111111111111111110011111111111100010001111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

	// top: 67, mid: 43, bot: 41
	reg[26799:0]top_text = 26800'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111011111111111111111111111110111111111111111111111111111111111111111111111111111111001111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111111111111111111101111111111111111111111111110011111011111111111111111111111111111111111111001101110111111111111101111111111111111111111111011111111111011111111111101111111111111111111111111111001111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111011111111111111111110111111111111111111111111111011111101111111111111111111111111111111111111111110111011111111111110111111111111111111111111101111111111101111111111110111111111111111111111111111101111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001101101110110000100011000001110001100001111100011000011100001000010000111000011100001100001000111010000000011000111000011111000001100001111000110110111000100001000011110000100001000011100001110000100001100011000010000110001110000111110000111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010010110111011001001101100110110110110011111101110110111111011100111111101100110110111110010011011101101110111011011011101111100110111111011011111010111011011011101111111101110011111110110011011011111011101101100111001110110110111011111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101011011101101110110110111011000001011111110111001011111101110111110000110111011001111011101101110110111011100000101110111110111011100001101111100111100000101110011111110111011111000011011101100111101110000010111101111000001011101111110000110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110001101110110111011011011101101111101111111011101101111110111011110111011011101111001101110110111011011101110111110111011111011101101110110111110101110111110111110011111011101111011101101110111100110111011111011110111101111101110111110111011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100110111011011101101100110110111110111111101110110111111011101111011001101110111110110111011011101101110111011111011101111100110110110011011111011011011111011111101111101110111101100110111011111011011101111101111011110111110111011111011001111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110011100001101110110110000011100011011111111000111011111110010111100000110111011000011011101101110111001100110001110000111110000111000001110001101100110001110010000111111001011110000011011101100001101111000110111101111100011100001111100000110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111110111111111101111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111011111111110111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111011101000010000011011101000011111000011000011000010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101101110110111001101101110110111111011101111110110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110010111011011101110110111011011111101110111000011011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011101101110111011011101101111110111011011101101110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101101110110111001101101110110111111011101101100110111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111000011100100001111000011100111110000110000011100100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011001111111111111111111111111111111111111111111111111111111111111111100110011111111111111111111111111111111111111111111111111111111111111111001100111111111111111111111111111111111111111111111111111111111111111100110011111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111110011001111111111111111110111111111111111111111111111111110000011111111100110011111111111111111000111111111111111111111111111111100000111111111001100111111111111111110001111111111111111111111111111110000011111111100110011111111111111111110111111111111111111111111111111100000011111111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111111011101111111111111111100011111111111111111111111111111111011101111111110111011111111111111111011001111111111111111111111111111110111011111111101110111111111111111110111011111111111111111111111111111011101111111110111011111111111111111110011111111111111111111111111111111110111111111101111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011101000000001100011000011111101111111111111111111111111111111101110110111010000000011000110000111111110111111111111111111111111111111011101101110100000000110001100001111111001111111111111111111111111111101110110111010000000011000110000111110101111111111111111111111111111111111011110001100001000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001101110110111011101101100111111110111111111111111111111111111111110000011011101101110111011011001111111110111111111111111111111111111111100000110111011011101110110110011111110001111111111111111111111111111110000011011101101110111011011001111111010111111111111111111111111111111111101110111011011111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111011011101110000010111111111011111111111111111111111111111111011101101110110111011100000101111111111011111111111111111111111111111110111011011101101110111000001011111111111011111111111111111111111111111011101101110110111011100000101111111011011111111111111111111111111111111110111011100101111000011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001011101101110111011111011111111101111111111111111111111111111111101110010111011011101110111110111111111011111111111111111111111111111111011100101110110111011101111101111111111101111111111111111111111111111101110010111011011101110111110111111100000011111111111111111111111111111111011101110110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101101110110111011101111101111111110111111111111111111111111111111110111011011101101110111011111011111110011111111111111111111111111111111101110110111011011101110111110111111101110111111111111111111111111111110111011011101101110111011111011111111110111111111111111111111111111111111101110111011011101100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111000011011101111000110111111100000111111111111111111111111111111000001110000110111011110001101111111000001111111111111111111111111111110000011100001101110111100011011111110000111111111111111111111111111111000001110000110111011110001101111111111011111111111111111111111111111111110111100011110010000011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[17199:0]mid_text = 17200'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111100111111111111111111111111111111111111111111111110111111111111111111111111101111111111111111111111111001111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101111111111111111111011111111111111111111111111100111111111111111111111111111100111111111111111111011111111111111111111111110111111111110111111111111001111111111111111111111111110000010000011110000111100111111011111111111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110111111111111111111101111111111111111111111111110111111111111111111111111111111111111111111111111101111111111111111111111111011111111111011111111111101111111111111111111111111111011111011101100111011110011111101111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011011011101100001000110000011100011000011111000110000111100001100011100011100011101001110110001110000111110000011000011110001101101110001000010000111100001000011000111000010001111101111101110010111111110101111110000011011101000000001100011100001110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110100101101110110010011011001101101101100111111011101101111110011101101101111101101110110110110110110111011111001101111110110111110101110110110111011111111011100111011101100100110111110000110111011011111111011011111001101101110110111011101110110011011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010110111011011101101101110110000010111111101110010111111011110000010111110000011011011011000001011101111101110111000011011111001111000001011100111111101110111101110010111011011111011111000011101100011101101111101110110111011011101110111001011101100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100011011101101110110110111011011111011111110111011011111101111011111011111011111101100101101111101110111110111011011101101111101011101111101111100111110111011110111011011101101111101111101111110111101100000011110111011011101101110111011101101110111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001101110110111011011001101101111101111111011101101111110111101111101111101111110111001110111110111011111001101101100110111110110110111110111111011111011101111011101101110110111110111110111111001110110111101111001101101110110111011101110110111011111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100111000011011101101101000111000110111111110001110111111011111000111000111000111011100111100011100001111100001110000011100011011001100011100100001111101110111110001110111011011111011111011111110000010011110111100000111000011100110011000111011101100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011001111111111111111111111111111111111111111111111111111111111111111100110011111111111111111111111111111111111111111111111111111111111111111001100111111111111111111111111111111111111111111111111111111111111111100110011111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111110011001111111111111111110111111111111111111111111111111110000011111111100110011111111111111111000111111111111111111111111111111100000111111111001100111111111111111110001111111111111111111111111111110000011111111100110011111111111111111110111111111111111111111111111111100000011111111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111111111011101111111111111111100011111111111111111111111111111111011101111111110111011111111111111111011001111111111111111111111111111110111011111111101110111111111111111110111011111111111111111111111111111011101111111110111011111111111111111110011111111111111111111111111111111110111111111101111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011101000000001100011000011111101111111111111111111111111111111101110110111010000000011000110000111111110111111111111111111111111111111011101101110100000000110001100001111111001111111111111111111111111111101110110111010000000011000110000111110101111111111111111111111111111111111011110001100001000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001101110110111011101101100111111110111111111111111111111111111111110000011011101101110111011011001111111110111111111111111111111111111111100000110111011011101110110110011111110001111111111111111111111111111110000011011101101110111011011001111111010111111111111111111111111111111111101110111011011111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111011011101110000010111111111011111111111111111111111111111111011101101110110111011100000101111111111011111111111111111111111111111110111011011101101110111000001011111111111011111111111111111111111111111011101101110110111011100000101111111011011111111111111111111111111111111110111011100101111000011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001011101101110111011111011111111101111111111111111111111111111111101110010111011011101110111110111111111011111111111111111111111111111111011100101110110111011101111101111111111101111111111111111111111111111101110010111011011101110111110111111100000011111111111111111111111111111111011101110110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101101110110111011101111101111111110111111111111111111111111111111110111011011101101110111011111011111110011111111111111111111111111111111101110110111011011101110111110111111101110111111111111111111111111111110111011011101101110111011111011111111110111111111111111111111111111111111101110111011011101100111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111000011011101111000110111111100000111111111111111111111111111111000001110000110111011110001101111111000001111111111111111111111111111110000011100001101110111100011011111110000111111111111111111111111111111000001110000110111011110001101111111111011111111111111111111111111111111110111100011110010000011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[16399:0]bot_text = 16400'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111001111111101111111111111111111111111111111111111101111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111011111111111111111110111111111111111111111111111001111111110111111111111111111111111111111111111110111111111111111111111111101111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101111111111111111111011111111111111111111111111101111111111011111111111111111111111111111111111111011111111111111111111111110111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110110111011000010001100000111000110000111110001100001111100001100001100011100000110000011100011100001111100000110000111100011011011100010000100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101001011011101100100110110011011011011001111110111011011111101110110011101110110011011001101101101101110111110011011111101101111101011101101101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110101101110110111011011011101100000101111111011100101111110111011011110111001011101101110110000010111011111011101110000110111110011110000010111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011000110111011011101101101110110111110111111101110110111111011101101111011101101110110111011011111011101111101110110111011011111010111011111011111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110011011101101110110110011011011111011111110111011011111101110110111101110110011011001101101111101110111110011011011001101111101101101111101111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111001110000110111011011000001110001101111111100011101111111000011011111000111000011100001111000111000011111000011100000111000110110011000111001000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111011111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011111111111111111111111111111111111111111111111111111111111111111001100111111111111111111111111111111111111111111111111111111111111111110011001111111111111111111111111111111111111111111111111111111111111111001100111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111100110011111111111111111101111111111111111111111111111111100000111111111001100111111111111111110001111111111111111111111111111111000001111111110011001111111111111111100011111111111111111111111111111100000111111111001100111111111111111111101111111111111111111111111111111000000111111110111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111110111011111111111111111000111111111111111111111111111111110111011111111101110111111111111111110110011111111111111111111111111111101110111111111011101111111111111111101110111111111111111111111111111110111011111111101110111111111111111111100111111111111111111111111111111111101111111111011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110110111010000000011000110000111111011111111111111111111111111111111011101101110100000000110001100001111111101111111111111111111111111111110111011011101000000001100011000011111110011111111111111111111111111111011101101110100000000110001100001111101011111111111111111111111111111111110111100011000010000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011011101101110111011011001111111101111111111111111111111111111111100000110111011011101110110110011111111101111111111111111111111111111111000001101110110111011101101100111111100011111111111111111111111111111100000110111011011101110110110011111110101111111111111111111111111111111111011101110110111111101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101101110110111011100000101111111110111111111111111111111111111111110111011011101101110111000001011111111110111111111111111111111111111111101110110111011011101110000010111111111110111111111111111111111111111110111011011101101110111000001011111110110111111111111111111111111111111111101110111001011110000111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110010111011011101110111110111111111011111111111111111111111111111111011100101110110111011101111101111111110111111111111111111111111111111110111001011101101110111011111011111111111011111111111111111111111111111011100101110110111011101111101111111000000111111111111111111111111111111110111011101101110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011011101101110111011111011111111101111111111111111111111111111111101110110111011011101110111110111111100111111111111111111111111111111111011101101110110111011101111101111111011101111111111111111111111111111101110110111011011101110111110111111111101111111111111111111111111111111111011101110110111011001110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110000110111011110001101111111000001111111111111111111111111111110000011100001101110111100011011111110000011111111111111111111111111111100000111000011011101111000110111111100001111111111111111111111111111110000011100001101110111100011011111111110111111111111111111111111111111111101111000111100100000111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	
	reg[2699:0]output_text = 2700'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111001111111111111111110011111100000111111111110011111111111111111111111111100111001111111111001111111111111111110011111100110011111111110011111111111111111111111111100111100100110010000010100011001100100000111100111001100001100001100001100111111111111111101111100100110011001110011001001100110011111100111001101100110011011100100111111111111111100111100100110011001110011001001100110011111100111001111100110011111100111111111111111111101111100100110011001110011001001100110011111100111001100000110011100000111111111111111111100111100100110011001110011001001100110011111100111001001100110011001100111111111111111111100111001100110011001110011001001100110011111100110011001100110011001000100111111111111111110000011110001011100010000011100000111001111100000111100000110001100000100111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[2699:0]input_text = 2700'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111001111110000001111111111001111111111111111111111111111111111111100111111111111111111111111001111110011100111111111001111111111111111111111111111111111111100110100011000001100111010000011110011100111000010000011000111001111111111111111111111111100110010011001100100111011001111110011110010110011001110110011001111111111111111111111111100110111011001100110111011001111110011110011110011001111110011111111111111111111111111111100110111001001100100111011001111110011110010000011001110000011111111111111111111111111111100110111001001100110111011001111110011100110010011001100110011111111111111111111111111111100110111001001100110110011001111110011100110110011001100110011001111111111111111111111111100110111001000001110001011100011110000001110000011100010000011001111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	reg[2796:0]buffer_text = 2797'b1111111111111111111111111111111111111111111111111111110011001111111111111111111111111111111111111111001100111111111111111111111111111111111111111100110011111111111111111111111111111111111111110011001111111111111111111111111111111111111111111111111111111111111111111100000111111111001100111111111111111111011111110000011111111100110011111111111111111000111111000001111111110011001111111111111111100011111100000111111111001100111111111111111111101111111111111111111111111111111111111111111111111011101111111110111011111111111111111000111111101110111111111011101111111111111111101100111110111011111111101110111111111111111110111011111011101111111110111011111111111111111110011111111111111111111111111111111111111111111111110111011011101000000001100011000011111101111111011101101110100000000110001100001111111101111101110110111010000000011000110000111111100111110111011011101000000001100011000011111010111111111111111111111111111111111111111111111111100000110111011011101110110110011111111011111110000011011101101110111011011001111111110111111000001101110110111011101101100111111100011111100000110111011011101110110110011111110101111111111111111111111111111111111111111111111111011101101110110111011100000101111111110111111101110110111011011101110000010111111111101111110111011011101101110111000001011111111111011111011101101110110111011100000101111111011011111111111111111111111111111111111111111111111110111001011101101110111011111011111111101111111011100101110110111011101111101111111110111111101110010111011011101110111110111111111110111110111001011101101110111011111011111110000001111111111111111111111111111111111111111111111101110110111011011101110111110111111111011111110111011011101101110111011111011111110011111111011101101110110111011101111101111111011101111101110110111011011101110111110111111111101111111111111111111111111111111111111111111111111000001110000110111011110001101111111000001111100000111000011011101111000110111111100000111110000011100001101110111100011011111110000111111000001110000110111011110001101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
	
	wire[15:0] H_counter;
	wire[15:0] V_counter;
	wire v_counter_trigger;
	
	assign hcount = H_counter + 144;
	assign vcount = V_counter + 35;
	
	horizontal_counter h_vga(clock_25, v_counter_trigger, H_counter);
	vertical_counter v_vga(clock_25, v_counter_trigger, V_counter);
	
	assign hsync = (H_counter > (640 + 15) && (H_counter < (640 + 16 + 95)));
	assign vsync = (V_counter > (480 + 9) && (V_counter < (480 + 10 + 1)));
	assign nsync = 1;
	
	assign red_sig = (hcount > 144 && hcount <= 783 && vcount > 35 && vcount <= 514) ? red : 0;
	assign green_sig = (hcount > 144 && hcount <= 783 && vcount > 35 && vcount <= 514) ? green : 0;
	assign blue_sig = (hcount > 144 && hcount <= 783 && vcount > 35 && vcount <= 514) ? blue : 0;
	
	always @(posedge clock_50) begin
		int_output_count1 = output_count1;
		int_output_count2 = output_count2;
		int_output_count3 = output_count3;
		int_output_count4 = output_count4;
		int_output_count_total = output_count1 + output_count2 + output_count3 + output_count4;
		int_received_count1 = received1;
		int_received_count2 = received2;
		int_received_count3 = received3;
		int_received_count4 = received4;
		int_received_count_total = int_received_count1 + int_received_count2 + int_received_count3 + int_received_count4;
		int_dropped_count1 = dropped1;
		int_dropped_count2 = dropped2;
		int_dropped_count3 = dropped3;
		int_dropped_count4 = dropped4;
		int_dropped_count_total = int_dropped_count1 + int_dropped_count2 + int_dropped_count3 + int_dropped_count4;
		
		if((hcount > 0+144) && (hcount <= 215+144+1+(383-360))) begin					    // LEFT BOX
			
			if((vcount > 0+35) && (vcount < 120+35)) begin 					 // INPUT BOX
				
				if((hcount > 30+144) && (hcount <= 120+144)) begin // INPUT TEXT
					if((vcount > 45+35) && (vcount <= 75+35)) begin
						red <= input_text[2699 - (90*(vcount-(46+35)) + (hcount-(31+144)))];
						green <= input_text[2699 - (90*(vcount-(46+35)) + (hcount-(31+144)))];
						blue <= input_text[2699 - (90*(vcount-(46+35)) + (hcount-(31+144)))];
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 120+144) && (hcount <= 140+144)) begin // INPUT DIG 3
					if((vcount > 45+35) && (vcount <= 75+35)) begin
						if(in_number[3] == 1) begin
							red <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(121+144)))];
							green <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(121+144)))];
							blue <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(121+144)))];
						end else if(in_number[3] == 0) begin
							red <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(121+144)))];
							green <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(121+144)))];
							blue <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(121+144)))];
						end else begin
							red <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(121+144)))];
							green <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(121+144)))];
							blue <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(121+144)))];
						end
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 140+144) && (hcount <= 160+144)) begin // INPUT DIG 2
					if((vcount > 45+35) && (vcount <= 75+35)) begin
						if(in_number[2] == 1) begin
							red <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(141+144)))];
							green <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(141+144)))];
							blue <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(141+144)))];
						end else if(in_number[2] == 0) begin
							red <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(141+144)))];
							green <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(141+144)))];
							blue <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(141+144)))];
						end else begin
							red <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(141+144)))];
							green <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(141+144)))];
							blue <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(141+144)))];
						end
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 160+144) && (hcount <= 180+144)) begin // INPUT DIG 1
					if((vcount > 45+35) && (vcount <= 75+35)) begin
						if(in_number[1] == 1) begin
							red <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(161+144)))];
							green <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(161+144)))];
							blue <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(161+144)))];
						end else if(in_number[1] == 0) begin
							red <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(161+144)))];
							green <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(161+144)))];
							blue <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(161+144)))];
						end else begin
							red <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(161+144)))];
							green <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(161+144)))];
							blue <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(161+144)))];
						end
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 180+144) && (hcount <= 200+144)) begin // INPUT DIG 0
					if((vcount > 45+35) && (vcount <= 75+35)) begin
						if(in_number[0] == 1) begin
							red <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(181+144)))];
							green <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(181+144)))];
							blue <= td_bir[599 - (20*(vcount-(46+35)) + (hcount-(181+144)))];
						end else if(in_number[0] == 0) begin
							red <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(181+144)))];
							green <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(181+144)))];
							blue <= td_sifir[599 - (20*(vcount-(46+35)) + (hcount-(181+144)))];
						end else begin
							red <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(181+144)))];
							green <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(181+144)))];
							blue <= td_dokuz[599 - (20*(vcount-(46+35)) + (hcount-(181+144)))];
						end
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else begin
					green <= 1;
					blue <= 1;
					red <= 1;
				end
			
			end else if((vcount >= 120+35) && (vcount <= 360+35+6)) begin 		 // BUFFERS BOX				
				
				if((hcount >= 40+144) && (hcount <= 80+144+1)) begin 				 // BUFFER 1 RED
					
					if((vcount > 35+120) && (vcount < 360+35+6) && hcount == 40+144) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if ((vcount > 35+120) && (vcount < 360+35+6) && hcount == 80+1+144) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 120+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 160+1+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 200+2+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					
					else if((vcount == 240+3+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 280+4+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 320+5+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 360+6+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount > 120+35) && (vcount <= 160+35)) begin 			 // DATA 1
						case(data1[17:15])
							3'b000: begin
								green <= 0;
								blue <= 0;
								red <= block_sifir[1599 - (40*(vcount-(121+35)) + (hcount-(41+144)))];
							end
							3'b001: begin
								green <= 0;
								blue <= 0;
								red <= block_bir[1599 - (40*(vcount-(121+35)) + (hcount-(41+144)))];
							end
							3'b010: begin
								green <= 0;
								blue <= 0;
								red <= block_iki[1599 - (40*(vcount-(121+35)) + (hcount-(41+144)))];
							end
							3'b011: begin
								green <= 0;
								blue <= 0;
								red <= block_uc[1599 - (40*(vcount-(121+35)) + (hcount-(41+144)))];
							end
							3'b100: begin
								green <= 1;
								blue <= 1;
								red <= 1;
							end
						endcase
					end else if((vcount > 160+35+1) && (vcount <= 200+35+1)) begin // DATA 2
						case(data1[14:12])
							3'b000: begin
								green <= 0;
								blue <= 0;
								red <= block_sifir[1599 - (40*(vcount-(161+35+1)) + (hcount-(41+144)))];
							end
							3'b001: begin
								green <= 0;
								blue <= 0;
								red <= block_bir[1599 - (40*(vcount-(161+35+1)) + (hcount-(41+144)))];
							end
							3'b010: begin
								green <= 0;
								blue <= 0;
								red <= block_iki[1599 - (40*(vcount-(161+35+1)) + (hcount-(41+144)))];
							end
							3'b011: begin
								green <= 0;
								blue <= 0;
								red <= block_uc[1599 - (40*(vcount-(161+35+1)) + (hcount-(41+144)))];
							end
							3'b100: begin
								green <= 1;
								blue <= 1;
								red <= 1;
							end
						endcase
					end else if((vcount > 200+35+2) && (vcount <= 240+35+2)) begin // DATA 3
						case(data1[11:9])
							3'b000: begin
								green <= 0;
								blue <= 0;
								red <= block_sifir[1599 - (40*(vcount-(201+35+2)) + (hcount-(41+144)))];
							end
							3'b001: begin
								green <= 0;
								blue <= 0;
								red <= block_bir[1599 - (40*(vcount-(201+35+2)) + (hcount-(41+144)))];
							end
							3'b010: begin
								green <= 0;
								blue <= 0;
								red <= block_iki[1599 - (40*(vcount-(201+35+2)) + (hcount-(41+144)))];
							end
							3'b011: begin
								green <= 0;
								blue <= 0;
								red <= block_uc[1599 - (40*(vcount-(201+35+2)) + (hcount-(41+144)))];
							end
							3'b100: begin
								green <= 1;
								blue <= 1;
								red <= 1;
							end
						endcase
					end else if((vcount > 240+35+3) && (vcount <= 280+35+3)) begin // DATA 4
						case(data1[8:6])
							3'b000: begin
								green <= 0;
								blue <= 0;
								red <= block_sifir[1599 - (40*(vcount-(241+35+3)) + (hcount-(41+144)))];
							end
							3'b001: begin
								green <= 0;
								blue <= 0;
								red <= block_bir[1599 - (40*(vcount-(241+35+3)) + (hcount-(41+144)))];
							end
							3'b010: begin
								green <= 0;
								blue <= 0;
								red <= block_iki[1599 - (40*(vcount-(241+35+3)) + (hcount-(41+144)))];
							end
							3'b011: begin
								green <= 0;
								blue <= 0;
								red <= block_uc[1599 - (40*(vcount-(241+35+3)) + (hcount-(41+144)))];
							end
							3'b100: begin
								green <= 1;
								blue <= 1;
								red <= 1;
							end
						endcase
					end else if((vcount > 280+35+4) && (vcount <= 320+35+4)) begin // DATA 5
						case(data1[5:3])
							3'b000: begin
								green <= 0;
								blue <= 0;
								red <= block_sifir[1599 - (40*(vcount-(281+35+4)) + (hcount-(41+144)))];
							end
							3'b001: begin
								green <= 0;
								blue <= 0;
								red <= block_bir[1599 - (40*(vcount-(281+35+4)) + (hcount-(41+144)))];
							end
							3'b010: begin
								green <= 0;
								blue <= 0;
								red <= block_iki[1599 - (40*(vcount-(281+35+4)) + (hcount-(41+144)))];
							end
							3'b011: begin
								green <= 0;
								blue <= 0;
								red <= block_uc[1599 - (40*(vcount-(281+35+4)) + (hcount-(41+144)))];
							end
							3'b100: begin
								green <= 1;
								blue <= 1;
								red <= 1;
							end
						endcase
					end else if((vcount > 320+35+5) && (vcount <= 360+35+5)) begin // DATA 6
						case(data1[2:0])
							3'b000: begin
								green <= 0;
								blue <= 0;
								red <= block_sifir[1599 - (40*(vcount-(321+35+5)) + (hcount-(41+144)))];
							end
							3'b001: begin
								green <= 0;
								blue <= 0;
								red <= block_bir[1599 - (40*(vcount-(321+35+5)) + (hcount-(41+144)))];
							end
							3'b010: begin
								green <= 0;
								blue <= 0;
								red <= block_iki[1599 - (40*(vcount-(321+35+5)) + (hcount-(41+144)))];
							end
							3'b011: begin
								green <= 0;
								blue <= 0;
								red <= block_uc[1599 - (40*(vcount-(321+35+5)) + (hcount-(41+144)))];
							end
							3'b100: begin
								green <= 1;
								blue <= 1;
								red <= 1;
							end
						endcase
					end
				
				end else if((hcount >= 85+144) && (hcount <= 125+144+1)) begin  // BUFFER 2 BLUE
				
				
				if((vcount > 35+120) && (vcount < 360+35+6) && hcount == 85+144) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if ((vcount > 35+120) && (vcount < 360+35+6) && hcount == 125+1+144) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 120+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 160+1+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 200+2+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					
					else if((vcount == 240+3+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 280+4+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 320+5+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 360+6+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					
					
				
					else if((vcount > 120+35) && (vcount <= 160+35)) begin 			 // DATA 1
						case(data2[17:15])
							3'b000: begin
								green <= 0;
								red <= 0;
								blue <= block_sifir[1599 - (40*(vcount-(121+35)) + (hcount-(86+144)))];
							end
							3'b001: begin
								green <= 0;
								red <= 0;
								blue <= block_bir[1599 - (40*(vcount-(121+35)) + (hcount-(86+144)))];
							end
							3'b010: begin
								green <= 0;
								red <= 0;
								blue <= block_iki[1599 - (40*(vcount-(121+35)) + (hcount-(86+144)))];
							end
							3'b011: begin
								green <= 0;
								red <= 0;
								blue <= block_uc[1599 - (40*(vcount-(121+35)) + (hcount-(86+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 160+35+1) && (vcount <= 200+35+1)) begin // DATA 2
						case(data2[14:12])
							3'b000: begin
								green <= 0;
								red <= 0;
								blue <= block_sifir[1599 - (40*(vcount-(161+35+1)) + (hcount-(86+144)))];
							end
							3'b001: begin
								green <= 0;
								red <= 0;
								blue <= block_bir[1599 - (40*(vcount-(161+35+1)) + (hcount-(86+144)))];
							end
							3'b010: begin
								green <= 0;
								red <= 0;
								blue <= block_iki[1599 - (40*(vcount-(161+35+1)) + (hcount-(86+144)))];
							end
							3'b011: begin
								green <= 0;
								red <= 0;
								blue <= block_uc[1599 - (40*(vcount-(161+35+1)) + (hcount-(86+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 200+35+2) && (vcount <= 240+35+2)) begin // DATA 3
						case(data2[11:9])
							3'b000: begin
								green <= 0;
								red <= 0;
								blue <= block_sifir[1599 - (40*(vcount-(201+35+2)) + (hcount-(86+144)))];
							end
							3'b001: begin
								green <= 0;
								red <= 0;
								blue <= block_bir[1599 - (40*(vcount-(201+35+2)) + (hcount-(86+144)))];
							end
							3'b010: begin
								green <= 0;
								red <= 0;
								blue <= block_iki[1599 - (40*(vcount-(201+35+2)) + (hcount-(86+144)))];
							end
							3'b011: begin
								green <= 0;
								red <= 0;
								blue <= block_uc[1599 - (40*(vcount-(201+35+2)) + (hcount-(86+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 240+35+3) && (vcount <= 280+35+3)) begin // DATA 4
						case(data2[8:6])
							3'b000: begin
								green <= 0;
								red <= 0;
								blue <= block_sifir[1599 - (40*(vcount-(241+35+3)) + (hcount-(86+144)))];
							end
							3'b001: begin
								green <= 0;
								red <= 0;
								blue <= block_bir[1599 - (40*(vcount-(241+35+3)) + (hcount-(86+144)))];
							end
							3'b010: begin
								green <= 0;
								red <= 0;
								blue <= block_iki[1599 - (40*(vcount-(241+35+3)) + (hcount-(86+144)))];
							end
							3'b011: begin
								green <= 0;
								red <= 0;
								blue <= block_uc[1599 - (40*(vcount-(241+35+3)) + (hcount-(86+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 280+35+4) && (vcount <= 320+35+4)) begin // DATA 5
						case(data2[5:3])
							3'b000: begin
								green <= 0;
								red <= 0;
								blue <= block_sifir[1599 - (40*(vcount-(281+35+4)) + (hcount-(86+144)))];
							end
							3'b001: begin
								green <= 0;
								red <= 0;
								blue <= block_bir[1599 - (40*(vcount-(281+35+4)) + (hcount-(86+144)))];
							end
							3'b010: begin
								green <= 0;
								red <= 0;
								blue <= block_iki[1599 - (40*(vcount-(281+35+4)) + (hcount-(86+144)))];
							end
							3'b011: begin
								green <= 0;
								red <= 0;
								blue <= block_uc[1599 - (40*(vcount-(281+35+4)) + (hcount-(86+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 320+35+5) && (vcount <= 360+35+5)) begin // DATA 6
						case(data2[2:0])
							3'b000: begin
								green <= 0;
								red <= 0;
								blue <= block_sifir[1599 - (40*(vcount-(321+35+5)) + (hcount-(86+144)))];
							end
							3'b001: begin
								green <= 0;
								red <= 0;
								blue <= block_bir[1599 - (40*(vcount-(321+35+5)) + (hcount-(86+144)))];
							end
							3'b010: begin
								green <= 0;
								red <= 0;
								blue <= block_iki[1599 - (40*(vcount-(321+35+5)) + (hcount-(86+144)))];
							end
							3'b011: begin
								green <= 0;
								red <= 0;
								blue <= block_uc[1599 - (40*(vcount-(321+35+5)) + (hcount-(86+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end
				
				end else if((hcount >= 130+144) && (hcount <= 170+144+1)) begin // BUFFER 3 YELLOW (RED + GREEN)
				
				if((vcount > 35+120) && (vcount < 360+35+6) && hcount == 130+144) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if ((vcount > 35+120) && (vcount < 360+35+6) && hcount == 170+1+144) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 120+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 160+1+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 200+2+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					
					else if((vcount == 240+3+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 280+4+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 320+5+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 360+6+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
			
					else if((vcount > 120+35) && (vcount <= 160+35)) begin 			 // DATA 1
						case(data3[17:15])
							3'b000: begin
								green <= block_sifir[1599 - (40*(vcount-(121+35)) + (hcount-(131+144)))];
								red <= block_sifir[1599 - (40*(vcount-(121+35)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b001: begin
								green <= block_bir[1599 - (40*(vcount-(121+35)) + (hcount-(131+144)))];
								red <= block_bir[1599 - (40*(vcount-(121+35)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b010: begin
								green <= block_iki[1599 - (40*(vcount-(121+35)) + (hcount-(131+144)))];
								red <= block_iki[1599 - (40*(vcount-(121+35)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b011: begin
								green <= block_uc[1599 - (40*(vcount-(121+35)) + (hcount-(131+144)))];
								red <= block_uc[1599 - (40*(vcount-(121+35)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 160+35+1) && (vcount <= 200+35+1)) begin // DATA 2
						case(data3[14:12])
							3'b000: begin
								green <= block_sifir[1599 - (40*(vcount-(161+35+1)) + (hcount-(131+144)))];
								red <= block_sifir[1599 - (40*(vcount-(161+35+1)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b001: begin
								green <= block_bir[1599 - (40*(vcount-(161+35+1)) + (hcount-(131+144)))];
								red <= block_bir[1599 - (40*(vcount-(161+35+1)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b010: begin
								green <= block_iki[1599 - (40*(vcount-(161+35+1)) + (hcount-(131+144)))];
								red <= block_iki[1599 - (40*(vcount-(161+35+1)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b011: begin
								green <= block_uc[1599 - (40*(vcount-(161+35+1)) + (hcount-(131+144)))];
								red <= block_uc[1599 - (40*(vcount-(161+35+1)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 200+35+2) && (vcount <= 240+35+2)) begin // DATA 3
						case(data3[11:9])
							3'b000: begin
								green <= block_sifir[1599 - (40*(vcount-(201+35+2)) + (hcount-(131+144)))];
								red <= block_sifir[1599 - (40*(vcount-(201+35+2)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b001: begin
								green <= block_bir[1599 - (40*(vcount-(201+35+2)) + (hcount-(131+144)))];
								red <= block_bir[1599 - (40*(vcount-(201+35+2)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b010: begin
								green <= block_iki[1599 - (40*(vcount-(201+35+2)) + (hcount-(131+144)))];
								red <= block_iki[1599 - (40*(vcount-(201+35+2)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b011: begin
								green <= block_uc[1599 - (40*(vcount-(201+35+2)) + (hcount-(131+144)))];
								red <= block_uc[1599 - (40*(vcount-(201+35+2)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 240+35+3) && (vcount <= 280+35+3)) begin // DATA 4
						case(data3[8:6])
							3'b000: begin
								green <= block_sifir[1599 - (40*(vcount-(241+35+3)) + (hcount-(131+144)))];
								red <= block_sifir[1599 - (40*(vcount-(241+35+3)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b001: begin
								green <= block_bir[1599 - (40*(vcount-(241+35+3)) + (hcount-(131+144)))];
								red <= block_bir[1599 - (40*(vcount-(241+35+3)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b010: begin
								green <= block_iki[1599 - (40*(vcount-(241+35+3)) + (hcount-(131+144)))];
								red <= block_iki[1599 - (40*(vcount-(241+35+3)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b011: begin
								green <= block_uc[1599 - (40*(vcount-(241+35+3)) + (hcount-(131+144)))];
								red <= block_uc[1599 - (40*(vcount-(241+35+3)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 280+35+4) && (vcount <= 320+35+4)) begin // DATA 5
						case(data3[5:3])
							3'b000: begin
								green <= block_sifir[1599 - (40*(vcount-(281+35+4)) + (hcount-(131+144)))];
								red <= block_sifir[1599 - (40*(vcount-(281+35+4)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b001: begin
								green <= block_bir[1599 - (40*(vcount-(281+35+4)) + (hcount-(131+144)))];
								red <= block_bir[1599 - (40*(vcount-(281+35+4)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b010: begin
								green <= block_iki[1599 - (40*(vcount-(281+35+4)) + (hcount-(131+144)))];
								red <= block_iki[1599 - (40*(vcount-(281+35+4)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b011: begin
								green <= block_uc[1599 - (40*(vcount-(281+35+4)) + (hcount-(131+144)))];
								red <= block_uc[1599 - (40*(vcount-(281+35+4)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 320+35+5) && (vcount <= 360+35+5)) begin // DATA 6
						case(data3[2:0])
							3'b000: begin
								green <= block_sifir[1599 - (40*(vcount-(321+35+5)) + (hcount-(131+144)))];
								red <= block_sifir[1599 - (40*(vcount-(321+35+5)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b001: begin
								green <= block_bir[1599 - (40*(vcount-(321+35+5)) + (hcount-(131+144)))];
								red <= block_bir[1599 - (40*(vcount-(321+35+5)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b010: begin
								green <= block_iki[1599 - (40*(vcount-(321+35+5)) + (hcount-(131+144)))];
								red <= block_iki[1599 - (40*(vcount-(321+35+5)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b011: begin
								green <= block_uc[1599 - (40*(vcount-(321+35+5)) + (hcount-(131+144)))];
								red <= block_uc[1599 - (40*(vcount-(321+35+5)) + (hcount-(131+144)))];
								blue <= 0;
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end
			
				end else if((hcount >= 175+144) && (hcount <= 215+144+1)) begin // BUFFER 4 GREEN
					if((vcount > 35+120) && (vcount < 360+35+6) && hcount == 175+144) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if ((vcount > 35+120) && (vcount < 360+35+6) && hcount == 215+1+144) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 120+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 160+1+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 200+2+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					
					else if((vcount == 240+3+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 280+4+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 320+5+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
					else if((vcount == 360+6+35)) begin
						green <= 0;
						blue <= 0;
						red <= 0;
					end
			
					else if((vcount > 120+35) && (vcount <= 160+35)) begin 			 // DATA 1
						case(data4[17:15])
							3'b000: begin
								blue <= 0;
								red <= 0;
								green <= block_sifir[1599 - (40*(vcount-(121+35)) + (hcount-(176+144)))];
							end
							3'b001: begin
								blue <= 0;
								red <= 0;
								green <= block_bir[1599 - (40*(vcount-(121+35)) + (hcount-(176+144)))];
							end
							3'b010: begin
								blue <= 0;
								red <= 0;
								green <= block_iki[1599 - (40*(vcount-(121+35)) + (hcount-(176+144)))];
							end
							3'b011: begin
								blue <= 0;
								red <= 0;
								green <= block_uc[1599 - (40*(vcount-(121+35)) + (hcount-(176+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 160+35+1) && (vcount <= 200+35+1)) begin // DATA 2
						case(data4[14:12])
							3'b000: begin
								blue <= 0;
								red <= 0;
								green <= block_sifir[1599 - (40*(vcount-(161+35+1)) + (hcount-(176+144)))];
							end
							3'b001: begin
								blue <= 0;
								red <= 0;
								green <= block_bir[1599 - (40*(vcount-(161+35+1)) + (hcount-(176+144)))];
							end
							3'b010: begin
								blue <= 0;
								red <= 0;
								green <= block_iki[1599 - (40*(vcount-(161+35+1)) + (hcount-(176+144)))];
							end
							3'b011: begin
								blue <= 0;
								red <= 0;
								green <= block_uc[1599 - (40*(vcount-(161+35+1)) + (hcount-(176+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 200+35+2) && (vcount <= 240+35+2)) begin // DATA 3
						case(data4[11:9])
							3'b000: begin
								blue <= 0;
								red <= 0;
								green <= block_sifir[1599 - (40*(vcount-(201+35+2)) + (hcount-(176+144)))];
							end
							3'b001: begin
								blue <= 0;
								red <= 0;
								green <= block_bir[1599 - (40*(vcount-(201+35+2)) + (hcount-(176+144)))];
							end
							3'b010: begin
								blue <= 0;
								red <= 0;
								green <= block_iki[1599 - (40*(vcount-(201+35+2)) + (hcount-(176+144)))];
							end
							3'b011: begin
								blue <= 0;
								red <= 0;
								green <= block_uc[1599 - (40*(vcount-(201+35+2)) + (hcount-(176+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 240+35+3) && (vcount <= 280+35+3)) begin // DATA 4
						case(data4[8:6])
							3'b000: begin
								blue <= 0;
								red <= 0;
								green <= block_sifir[1599 - (40*(vcount-(241+35+3)) + (hcount-(176+144)))];
							end
							3'b001: begin
								blue <= 0;
								red <= 0;
								green <= block_bir[1599 - (40*(vcount-(241+35+3)) + (hcount-(176+144)))];
							end
							3'b010: begin
								blue <= 0;
								red <= 0;
								green <= block_iki[1599 - (40*(vcount-(241+35+3)) + (hcount-(176+144)))];
							end
							3'b011: begin
								blue <= 0;
								red <= 0;
								green <= block_uc[1599 - (40*(vcount-(241+35+3)) + (hcount-(176+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 280+35+4) && (vcount <= 320+35+4)) begin // DATA 5
						case(data4[5:3])
							3'b000: begin
								blue <= 0;
								red <= 0;
								green <= block_sifir[1599 - (40*(vcount-(281+35+4)) + (hcount-(176+144)))];
							end
							3'b001: begin
								blue <= 0;
								red <= 0;
								green <= block_bir[1599 - (40*(vcount-(281+35+4)) + (hcount-(176+144)))];
							end
							3'b010: begin
								blue <= 0;
								red <= 0;
								green <= block_iki[1599 - (40*(vcount-(281+35+4)) + (hcount-(176+144)))];
							end
							3'b011: begin
								blue <= 0;
								red <= 0;
								green <= block_uc[1599 - (40*(vcount-(281+35+4)) + (hcount-(176+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end else if((vcount > 320+35+5) && (vcount <= 360+35+5)) begin // DATA 6
						case(data4[2:0])
							3'b000: begin
								blue <= 0;
								red <= 0;
								green <= block_sifir[1599 - (40*(vcount-(321+35+5)) + (hcount-(176+144)))];
							end
							3'b001: begin
								blue <= 0;
								red <= 0;
								green <= block_bir[1599 - (40*(vcount-(321+35+5)) + (hcount-(176+144)))];
							end
							3'b010: begin
								blue <= 0;
								red <= 0;
								green <= block_iki[1599 - (40*(vcount-(321+35+5)) + (hcount-(176+144)))];
							end
							3'b011: begin
								blue <= 0;
								red <= 0;
								green <= block_uc[1599 - (40*(vcount-(321+35+5)) + (hcount-(176+144)))];
							end
							3'b100: begin
								green <= 1;
								red <= 1;
								blue <= 1;
							end
						endcase
					end
			
				end else begin // SPACE BTW BUFFERS
					red <= 1;
					green <= 1;
					blue <= 1;
				end
			end else if ((vcount >= 360+35+5) && (vcount <= 371+35+5+5)) begin
				if((hcount > 144) && (hcount <= 227+144)) begin // buffer text 
					if((vcount > 360+35+5+5) && (vcount <= 360+35+5+5+11)) begin
						red <= buffer_text[2496 - (227*(vcount-(370+35+1)) + (hcount-(1+144)))];
						green <= buffer_text[2496 - (227*(vcount-(370+35+1)) + (hcount-(1+144)))];
						blue <= buffer_text[2496 - (227*(vcount-(370+35+1)) + (hcount-(1+144)))];
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end
			
			end else if((vcount > 371+35+5+5) && (vcount <= 480+35)) begin // OUTPUT BOX
								
				if((hcount > 30+144) && (hcount <= 120+144)) begin // OUTPUT TEXT
					if((vcount > 405+35) && (vcount <= 435+35)) begin
						red <= output_text[2699 - (90*(vcount-(406+35)) + (hcount-(31+144)))];
						green <= output_text[2699 - (90*(vcount-(406+35)) + (hcount-(31+144)))];
						blue <= output_text[2699 - (90*(vcount-(406+35)) + (hcount-(31+144)))];
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 120+144) && (hcount <= 140+144)) begin // OUTPUT DIG 3
					if((vcount > 405+35) && (vcount <= 435+35)) begin
						if(outputted_buffer_packet[3] == 1) begin
							red <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(121+144)))];
							green <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(121+144)))];
							blue <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(121+144)))];
						end else if(outputted_buffer_packet[3] == 0) begin
							red <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(121+144)))];
							green <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(121+144)))];
							blue <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(121+144)))];
						end else begin
							red <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(121+144)))];
							green <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(121+144)))];
							blue <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(121+144)))];
						end
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 140+144) && (hcount <= 160+144)) begin // OUTPUT DIG 2
					if((vcount > 405+35) && (vcount <= 435+35)) begin
						if(outputted_buffer_packet[2] == 1) begin
							red <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(141+144)))];
							green <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(141+144)))];
							blue <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(141+144)))];
						end else if(outputted_buffer_packet[2] == 0) begin
							red <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(141+144)))];
							green <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(141+144)))];
							blue <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(141+144)))];
						end else begin
							red <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(141+144)))];
							green <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(141+144)))];
							blue <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(141+144)))];
						end
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 160+144) && (hcount <= 180+144)) begin // OUTPUT DIG 1
					if((vcount > 405+35) && (vcount <= 435+35)) begin
						if(outputted_buffer_packet[1] == 1) begin
							red <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(161+144)))];
							green <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(161+144)))];
							blue <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(161+144)))];
						end else if(outputted_buffer_packet[1] == 0) begin
							red <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(161+144)))];
							green <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(161+144)))];
							blue <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(161+144)))];
						end else begin
							red <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(161+144)))];
							green <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(161+144)))];
							blue <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(161+144)))];
						end
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 180+144) && (hcount <= 200+144)) begin // OUTPUT DIG 0
					if((vcount > 405+35) && (vcount <= 435+35)) begin
						if(outputted_buffer_packet[0] == 1) begin
							red <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(181+144)))];
							green <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(181+144)))];
							blue <= td_bir[599 - (20*(vcount-(406+35)) + (hcount-(181+144)))];
						end else if(outputted_buffer_packet[0] == 0) begin
							red <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(181+144)))];
							green <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(181+144)))];
							blue <= td_sifir[599 - (20*(vcount-(406+35)) + (hcount-(181+144)))];
						end else begin
							red <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(181+144)))];
							green <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(181+144)))];
							blue <= td_dokuz[599 - (20*(vcount-(406+35)) + (hcount-(181+144)))];
						end
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else begin
					green <= 1;
					blue <= 1;
					red <= 1;
				end
				
			end else begin
				green <= 1;
				blue <= 1;
				red <= 1;
			end
			
		end else if((hcount > 239+144) && (hcount <= 640+144)) begin // RIGHT BOX
			
			if((vcount > 28+35) && (vcount <= 95+35)) begin // TOP TEXT
			
				red <= top_text[26799 - (400*(vcount-(29+35)) + (hcount-(240+144)))];
				green <= top_text[26799 - (400*(vcount-(29+35)) + (hcount-(240+144)))];
				blue <= top_text[26799 - (400*(vcount-(29+35)) + (hcount-(240+144)))];
				
			end else if((vcount > 95+35) && (vcount <= 125+35)) begin // TOP DIGS
			
				if((hcount > 270+144) && (hcount <= 330+144)) begin // output_count1
					if((hcount > 270+144) && (hcount <= 290+144)) begin // output_count1 dig 2
						dumdig = int_output_count1 / 100;
						case(dumdig)
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(271+144)))];
							end
						endcase
					end else if((hcount > 290+144) && (hcount <= 310+144)) begin // output_count1 dig 1
						dumdig = (int_output_count1 - 100*(int_output_count1 / 100))/10;
						case(dumdig)
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(291+144)))];
							end
						endcase
					end else if((hcount > 310+144) && (hcount <= 330+144)) begin // output_count1 dig 0
						dumdig = int_output_count1 - 10*(int_output_count1/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(311+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 341+144) && (hcount <= 401+144)) begin // output_count2
					if((hcount > 341+144) && (hcount <= 361+144)) begin // output_count2 dig 2
						dumdig = int_output_count2 / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(342+144)))];
							end
						endcase
					end else if((hcount > 361+144) && (hcount <= 381+144)) begin // output_count2 dig 1
						dumdig = (int_output_count2 - 100*(int_output_count2 / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(362+144)))];
							end
						endcase
					end else if((hcount > 381+144) && (hcount <= 401+144)) begin // output_count2 dig 0
						dumdig = int_output_count2 - 10*(int_output_count2/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(382+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 412+144) && (hcount <= 472+144)) begin // output_count3
					if((hcount > 412+144) && (hcount <= 432+144)) begin // output_count3 dig 2
						dumdig = int_output_count3 / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(413+144)))];
							end
						endcase
					end else if((hcount > 432+144) && (hcount <= 452+144)) begin // output_count3 dig 1
						dumdig = (int_output_count3 - 100*(int_output_count3 / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(433+144)))];
							end
						endcase
					end else if((hcount > 452+144) && (hcount <= 472+144)) begin // output_count3 dig 0
						dumdig = int_output_count3 - 10*(int_output_count3/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(453+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 482+144) && (hcount <= 542+144)) begin // output_count4
					if((hcount > 482+144) && (hcount <= 502+144)) begin // output_count4 dig 2
						dumdig = int_output_count4 / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(483+144)))];
							end
						endcase
					end else if((hcount > 502+144) && (hcount <= 522+144)) begin // output_count4 dig 1
						dumdig = (int_output_count4 - 100*(int_output_count4 / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(503+144)))];
							end
						endcase
					end else if((hcount > 522+144) && (hcount <= 542+144)) begin // output_count4 dig 0
						dumdig = int_output_count4 - 10*(int_output_count4/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(523+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 554+144) && (hcount <= 614+144)) begin // output_count_total
					if((hcount > 554+144) && (hcount <= 574+144)) begin // output_count_total dig 2
						dumdig = int_output_count_total / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(555+144)))];
							end
						endcase
					end else if((hcount > 574+144) && (hcount <= 594+144)) begin // output_count_total dig 1
						dumdig = (int_output_count_total - 100*(int_output_count_total / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(575+144)))];
							end
						endcase
					end else if((hcount > 594+144) && (hcount <= 614+144)) begin // output_count_total dig 0
						dumdig = int_output_count_total - 10*(int_output_count_total/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_sifir[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_bir[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_iki[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_uc[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_dort[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_bes[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_alti[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_yedi[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_sekiz[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								green <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
								blue <= td_dokuz[599 - (20*(vcount-(96+35)) + (hcount-(595+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else begin
					green <= 1;
					blue <= 1;
					red <= 1;
				end
			end else if((vcount > 194+35) && (vcount <= 237+35)) begin // MID TEXT
			
				red <= mid_text[17199 - (400*(vcount-(195+35)) + (hcount-(240+144)))];
				green <= mid_text[17199 - (400*(vcount-(195+35)) + (hcount-(240+144)))];
				blue <= mid_text[17199 - (400*(vcount-(195+35)) + (hcount-(240+144)))];
			
			end else if((vcount > 237+35) && (vcount <= 267+35)) begin // MID DIGS
			
				if((hcount > 270+144) && (hcount <= 330+144)) begin // received_count1
					if((hcount > 270+144) && (hcount <= 290+144)) begin // received_count1 dig 2
						dumdig = int_received_count1 / 100;
						case(dumdig)
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(271+144)))];
							end
						endcase
					end else if((hcount > 290+144) && (hcount <= 310+144)) begin // received_count1 dig 1
						dumdig = (int_received_count1 - 100*(int_received_count1 / 100))/10;
						case(dumdig)
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(291+144)))];
							end
						endcase
					end else if((hcount > 310+144) && (hcount <= 330+144)) begin // received_count1 dig 0
						dumdig = int_received_count1 - 10*(int_received_count1/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(311+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 341+144) && (hcount <= 401+144)) begin // received_count2
					if((hcount > 341+144) && (hcount <= 361+144)) begin // received_count2 dig 2
						dumdig = int_received_count2 / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(342+144)))];
							end
						endcase
					end else if((hcount > 361+144) && (hcount <= 381+144)) begin // received_count2 dig 1
						dumdig = (int_received_count2 - 100*(int_received_count2 / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(362+144)))];
							end
						endcase
					end else if((hcount > 381+144) && (hcount <= 401+144)) begin // received_count2 dig 0
						dumdig = int_received_count2 - 10*(int_received_count2/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(382+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 412+144) && (hcount <= 472+144)) begin // received_count3
					if((hcount > 412+144) && (hcount <= 432+144)) begin // received_count3 dig 2
						dumdig = int_received_count3 / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(413+144)))];
							end
						endcase
					end else if((hcount > 432+144) && (hcount <= 452+144)) begin // received_count3 dig 1
						dumdig = (int_received_count3 - 100*(int_received_count3 / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(433+144)))];
							end
						endcase
					end else if((hcount > 452+144) && (hcount <= 472+144)) begin // received_count3 dig 0
						dumdig = int_received_count3 - 10*(int_received_count3/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(453+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 482+144) && (hcount <= 542+144)) begin // received_count4
					if((hcount > 482+144) && (hcount <= 502+144)) begin // received_count4 dig 2
						dumdig = int_received_count4 / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(483+144)))];
							end
						endcase
					end else if((hcount > 502+144) && (hcount <= 522+144)) begin // received_count4 dig 1
						dumdig = (int_received_count4 - 100*(int_received_count4 / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(503+144)))];
							end
						endcase
					end else if((hcount > 522+144) && (hcount <= 542+144)) begin // received_count4 dig 0
						dumdig = int_received_count4 - 10*(int_received_count4/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(523+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 554+144) && (hcount <= 614+144)) begin // received_count_total
					if((hcount > 554+144) && (hcount <= 574+144)) begin // received_count_total dig 2
						dumdig = int_received_count_total / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(555+144)))];
							end
						endcase
					end else if((hcount > 574+144) && (hcount <= 594+144)) begin // received_count_total dig 1
						dumdig = (int_received_count_total - 100*(int_received_count_total / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(575+144)))];
							end
						endcase
					end else if((hcount > 594+144) && (hcount <= 614+144)) begin // received_count_total dig 0
						dumdig = int_received_count_total - 10*(int_received_count_total/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_sifir[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_bir[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_iki[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_uc[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_dort[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_bes[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_alti[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_yedi[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 142-(96+35)) + (hcount-(595+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else begin
					green <= 1;
					blue <= 1;
					red <= 1;
				end
				
			end else if((vcount > 333+35) && (vcount <= 374+35)) begin // BOT TEXT
			
				red <= bot_text[16399 - (400*(vcount-(334+35)) + (hcount-(240+144)))];
				green <= bot_text[16399 - (400*(vcount-(334+35)) + (hcount-(240+144)))];
				blue <= bot_text[16399 - (400*(vcount-(334+35)) + (hcount-(240+144)))];
			
			end else if((vcount > 374+35) && (vcount <= 404+35)) begin // BOT DIGS
				
				if((hcount > 270+144) && (hcount <= 330+144)) begin // dropped_count1
					if((hcount > 270+144) && (hcount <= 290+144)) begin // dropped_count1 dig 2
						dumdig = int_dropped_count1 / 100;
						case(dumdig)
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(271+144)))];
							end
						endcase
					end else if((hcount > 290+144) && (hcount <= 310+144)) begin // dropped_count1 dig 1
						dumdig = (int_dropped_count1 - 100*(int_dropped_count1 / 100))/10;
						case(dumdig)
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(291+144)))];
							end
						endcase
					end else if((hcount > 310+144) && (hcount <= 330+144)) begin // dropped_count1 dig 0
						dumdig = int_dropped_count1 - 10*(int_dropped_count1/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(311+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 341+144) && (hcount <= 401+144)) begin // dropped_count2
					if((hcount > 341+144) && (hcount <= 361+144)) begin // dropped_count2 dig 2
						dumdig = int_dropped_count2 / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(342+144)))];
							end
						endcase
					end else if((hcount > 361+144) && (hcount <= 381+144)) begin // dropped_count2 dig 1
						dumdig = (int_dropped_count2 - 100*(int_dropped_count2 / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(362+144)))];
							end
						endcase
					end else if((hcount > 381+144) && (hcount <= 401+144)) begin // dropped_count2 dig 0
						dumdig = int_dropped_count2 - 10*(int_dropped_count2/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(382+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 412+144) && (hcount <= 472+144)) begin // dropped_count3
					if((hcount > 412+144) && (hcount <= 432+144)) begin // dropped_count3 dig 2
						dumdig = int_dropped_count3 / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(413+144)))];
							end
						endcase
					end else if((hcount > 432+144) && (hcount <= 452+144)) begin // dropped_count3 dig 1
						dumdig = (int_dropped_count3 - 100*(int_dropped_count3 / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(433+144)))];
							end
						endcase
					end else if((hcount > 452+144) && (hcount <= 472+144)) begin // dropped_count3 dig 0
						dumdig = int_dropped_count3 - 10*(int_dropped_count3/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(453+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 482+144) && (hcount <= 542+144)) begin // dropped_count4
					if((hcount > 482+144) && (hcount <= 502+144)) begin // dropped_count4 dig 2
						dumdig = int_dropped_count4 / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(483+144)))];
							end
						endcase
					end else if((hcount > 502+144) && (hcount <= 522+144)) begin // dropped_count4 dig 1
						dumdig = (int_dropped_count4 - 100*(int_dropped_count4 / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(503+144)))];
							end
						endcase
					end else if((hcount > 522+144) && (hcount <= 542+144)) begin // dropped_count4 dig 0
						dumdig = int_dropped_count4 - 10*(int_dropped_count4/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(523+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else if((hcount > 554+144) && (hcount <= 614+144)) begin // dropped_count_total
					if((hcount > 554+144) && (hcount <= 574+144)) begin // dropped_count_total dig 2
						dumdig = int_dropped_count_total / 100;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(555+144)))];
							end
						endcase
					end else if((hcount > 574+144) && (hcount <= 594+144)) begin // dropped_count_total dig 1
						dumdig = (int_dropped_count_total - 100*(int_dropped_count_total / 100))/10;
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(575+144)))];
							end
						endcase
					end else if((hcount > 594+144) && (hcount <= 614+144)) begin // dropped_count_total dig 0
						dumdig = int_dropped_count_total - 10*(int_dropped_count_total/10);
						case(dumdig) 
							0: begin
								red <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_sifir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
							1: begin
								red <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_bir[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
							2: begin
								red <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_iki[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
							3: begin
								red <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_uc[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
							4: begin
								red <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_dort[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
							5: begin
								red <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_bes[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
							6: begin
								red <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_alti[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
							7: begin
								red <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_yedi[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
							8: begin
								red <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_sekiz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
							9: begin
								red <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								green <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
								blue <= td_dokuz[599 - (20*(vcount - 137 - 142-(96+35)) + (hcount-(595+144)))];
							end
						endcase
					end else begin
						green <= 1;
						blue <= 1;
						red <= 1;
					end
				end else begin
					green <= 1;
					blue <= 1;
					red <= 1;
				end
				
			end else begin
				red <= 1;
				green <= 1;
				blue <= 1;
			end
			
		end
		
	end
	
endmodule
